module NameSuite_InputPortNameComp_1(
    input [19:0] io_in,
    output[19:0] io_out
);


  assign io_out = io_in;
endmodule

