module ZeroWidthTest_ZeroWidthForceMatching_1(
    output io
);



  assign io = 1'h0;
endmodule

