module NameSuite_BindFourthComp_1(
    input [4:0] io_in,
    output [4:0] io_out
);


  assign io_out = io_in;
endmodule

